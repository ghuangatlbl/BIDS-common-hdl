//https://forums.xilinx.com/t5/Welcome-Join/synthesizable-verilog-connecting-inout-pins/td-p/284628
module via (.a(w), .b(w));
inout w;
wire w;
endmodule
